library ieee;
use ieee.std_logic_1164.all;
use ieee.math_real.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity Top_Module is
	port (
		clk : in std_logic;
		rst : in std_logic;
	);
end entity;

architecture behavioral of Top_Module is

begin
	Top_ModuleInst : process (clk)
	begin
		if rising_edge(clk) then
		end if;
	end process; -- Top_ModuleInst
end architecture;
